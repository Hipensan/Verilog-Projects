library verilog;
use verilog.vl_types.all;
entity tb_segment is
end tb_segment;
