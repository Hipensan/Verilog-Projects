module (
	input
	output
	);


// params



// nets



// regs



// subModules




// FSM







endmodule